library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.fixed_float_types.all; -- package virgule fixe
use ieee.fixed_pkg.all;
use ieee.math_real.all;         -- bibliothèque mathématique pour la trigonométrie
use work.types.all;             -- types prédéfinis

entity testbench is
end entity testbench;
